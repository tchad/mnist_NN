/*
"""
    EE278: Miniproject 4, RTL Implementation of the Inference Engine
           for MNIST Digit Recognition 
    SJSU, Fall 2018
    Tomasz Chadzynski
"""
*/


package util_fix;
    enum { SCALER_DIV, SCALER_MUL } scaler_t;
endpackage
